------------------------------------------------------------------------------------
---- Company: 
---- Engineer: 
---- 
---- Create Date:    18:29:29 03/31/2018 
---- Design Name: 
---- Module Name:    data_input - Behavioral 
---- Project Name: 	 
---- Target Devices: 
---- Tool versions: 
---- Description: 
----
---- Dependencies: 
----
---- Revision: 
---- Revision 0.01 - File Created
---- Additional Comments: 
----
------------------------------------------------------------------------------------
--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--
---- Uncomment the following library declaration if using
---- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;
--
---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
----library UNISIM;
----use UNISIM.VComponents.all;
--
--entity data_input is
--    Port ( serial_clock : in  STD_LOGIC;
--           serial_data : in  STD_LOGIC;
--           reset : in  STD_LOGIC;
--           full_byte : out  STD_LOGIC;
--           data_recv : out  STD_LOGIC_VECTOR (7 downto 0));
--end data_input;
--
--architecture Behavioral of data_input is
--
--	signal reg : std_logic_vector( 7 downto 0 );
--	signal ctr : unsigned( 2 downto 0 );
--
--begin
--
--	data_recv <= reg;
--	full_byte <= '1' when ctr = 7 else '0';
--
--	shifter : process( serial_clock, reset ) 
--	begin
--		
--		if( reset = '1' ) then
--			ctr <= 0;
--			reg <= ( others => '0' );
--			
--		elsif( serial_clock'event and serial_clock = '1' ) then
--			
--			if( ctr < 7 ) then
--				reg <= reg( 46 downto 0 ) & serial_data;
--				ctr <= ctr +1;
--			end if;
--			
--		end if;
--		
--	end process shifter;
--
--end Behavioral;
--
